`timescale 1 ps / 1 ps
`define RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE_REG_INIT
`define RANDOMIZE_DELAY 10
/*
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
*/

module simulation_top
(
    
);
reg    cpu_clk;
reg    cpu_reset;
wire    ddr4_init_copmlete;
wire    flash_int;
wire    uart_int;

	initial begin
		cpu_clk = 1'b0;
		cpu_reset = 1'b1;
		# 777.7
		cpu_reset = 1'b0;

		//# 2000000
		//$finish;
	end

  always begin
		#(10) cpu_clk = ~cpu_clk;
	end

  assign ddr4_init_copmlete = 1'b1;
  assign flash_int = 1'b0;
  assign uart_int = 1'b0;

wire           mem_axi_1_aw_ready;
assign    mem_axi_1_aw_ready = 'd1;
wire           mem_axi_1_aw_valid;
wire    [3:0]  mem_axi_1_aw_bits_id;
wire    [35:0] mem_axi_1_aw_bits_addr;
wire    [7:0]  mem_axi_1_aw_bits_len;
wire    [2:0]  mem_axi_1_aw_bits_size;
wire    [1:0]  mem_axi_1_aw_bits_burst;
wire           mem_axi_1_aw_bits_lock;
wire    [3:0]  mem_axi_1_aw_bits_cache;
wire    [2:0]  mem_axi_1_aw_bits_prot;
wire    [3:0]  mem_axi_1_aw_bits_qos;
wire           mem_axi_1_w_ready;
assign    mem_axi_1_w_ready = 'd1;
wire           mem_axi_1_w_valid;
wire    [63:0] mem_axi_1_w_bits_data;
wire    [7:0]  mem_axi_1_w_bits_strb;
wire           mem_axi_1_w_bits_last;
wire           mem_axi_1_b_ready;
wire           mem_axi_1_b_valid;
wire    [3:0]  mem_axi_1_b_bits_id;
wire    [1:0]  mem_axi_1_b_bits_resp;
assign    mem_axi_1_b_valid = 'd0;
assign    mem_axi_1_b_bits_id = 'd0;
assign    mem_axi_1_b_bits_resp = 'd0;
wire           mem_axi_1_ar_ready;
assign    mem_axi_1_ar_ready = 'd1;
wire           mem_axi_1_ar_valid;
wire    [3:0]  mem_axi_1_ar_bits_id;
wire    [35:0] mem_axi_1_ar_bits_addr;
wire    [7:0]  mem_axi_1_ar_bits_len;
wire    [2:0]  mem_axi_1_ar_bits_size;
wire    [1:0]  mem_axi_1_ar_bits_burst;
wire           mem_axi_1_ar_bits_lock;
wire    [3:0]  mem_axi_1_ar_bits_cache;
wire    [2:0]  mem_axi_1_ar_bits_prot;
wire    [3:0]  mem_axi_1_ar_bits_qos;
wire           mem_axi_1_r_ready;
wire           mem_axi_1_r_valid;
wire    [3:0]  mem_axi_1_r_bits_id;
wire    [63:0] mem_axi_1_r_bits_data;
wire    [1:0]  mem_axi_1_r_bits_resp;
wire           mem_axi_1_r_bits_last;
assign    mem_axi_1_r_valid = 'd0;
assign    mem_axi_1_r_bits_id = 'd0;
assign    mem_axi_1_r_bits_data = 'd0;
assign    mem_axi_1_r_bits_resp = 'd0;
assign    mem_axi_1_r_bits_last = 'd0;

wire           mmio_axi_0_aw_ready;
assign    mmio_axi_0_aw_ready = 'd1;
wire           mmio_axi_0_aw_valid;
wire    [3:0]  mmio_axi_0_aw_bits_id;
wire    [31:0] mmio_axi_0_aw_bits_addr;
wire    [7:0]  mmio_axi_0_aw_bits_len;
wire    [2:0]  mmio_axi_0_aw_bits_size;
wire    [1:0]  mmio_axi_0_aw_bits_burst;
wire           mmio_axi_0_aw_bits_lock;
wire    [3:0]  mmio_axi_0_aw_bits_cache;
wire    [2:0]  mmio_axi_0_aw_bits_prot;
wire    [3:0]  mmio_axi_0_aw_bits_qos;
wire           mmio_axi_0_w_ready;
assign    mmio_axi_0_w_ready = 'd1;
wire           mmio_axi_0_w_valid;
wire    [63:0] mmio_axi_0_w_bits_data;
wire    [7:0]  mmio_axi_0_w_bits_strb;
wire           mmio_axi_0_w_bits_last;
wire           mmio_axi_0_b_ready;
wire           mmio_axi_0_b_valid;
wire    [3:0]  mmio_axi_0_b_bits_id;
wire    [1:0]  mmio_axi_0_b_bits_resp;
assign    mmio_axi_0_b_bits_id = 'd0;
assign    mmio_axi_0_b_valid = 'd0;
assign    mmio_axi_0_b_bits_resp = 'd0;
wire           mmio_axi_0_ar_ready;
assign    mmio_axi_0_ar_ready = 'd1;
wire           mmio_axi_0_ar_valid;
wire    [3:0]  mmio_axi_0_ar_bits_id;
wire    [31:0] mmio_axi_0_ar_bits_addr;
wire    [7:0]  mmio_axi_0_ar_bits_len;
wire    [2:0]  mmio_axi_0_ar_bits_size;
wire    [1:0]  mmio_axi_0_ar_bits_burst;
wire           mmio_axi_0_ar_bits_lock;
wire    [3:0]  mmio_axi_0_ar_bits_cache;
wire    [2:0]  mmio_axi_0_ar_bits_prot;
wire    [3:0]  mmio_axi_0_ar_bits_qos;
wire           mmio_axi_0_r_ready;
wire           mmio_axi_0_r_valid;
wire    [3:0]  mmio_axi_0_r_bits_id;
wire    [63:0] mmio_axi_0_r_bits_data;
wire    [1:0]  mmio_axi_0_r_bits_resp;
wire           mmio_axi_0_r_bits_last;
assign    mmio_axi_0_r_valid = 'd0;
assign    mmio_axi_0_r_bits_id = 'd0;
assign    mmio_axi_0_r_bits_data = 'd0;
assign    mmio_axi_0_r_bits_resp = 'd0;
assign    mmio_axi_0_r_bits_last = 'd0;

SERVETop SERVETop(
  .clock (cpu_clk), // @[:freedom.serve.SERVEiFPGAConfig.fir@561594.4]
  .reset (cpu_reset | ~ddr4_init_copmlete), // @[:freedom.serve.SERVEiFPGAConfig.fir@561595.4]
  /*. io_ps_axi_slave_aw_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_aw_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_aw_bits_id ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_aw_bits_addr ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_aw_bits_len ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_aw_bits_size ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_aw_bits_burst ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_aw_bits_lock ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_aw_bits_cache ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_aw_bits_prot ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_aw_bits_qos ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_w_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_w_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_w_bits_data ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_w_bits_strb ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_w_bits_last ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_b_ready (1'b1), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_b_valid (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_b_bits_id (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_b_bits_resp (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_ar_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_ar_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_ar_bits_id ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_ar_bits_addr ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_ar_bits_len ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_ar_bits_size ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_ar_bits_burst ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_ar_bits_lock ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_ar_bits_cache ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_ar_bits_prot ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_ar_bits_qos ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_r_ready ('d1), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_r_valid (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_r_bits_id (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_r_bits_data (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_r_bits_resp (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_ps_axi_slave_r_bits_last (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]*/
  .io_mac_int ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_sdio_int ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_uart_int (uart_int), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .io_usb_int ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  //.io_jtag_TCK ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  //.io_jtag_TMS ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  //.io_jtag_TDI ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  //.io_jtag_TDO_data ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  //.io_jtag_TDO_driven ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  //.io_gpio_btns ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  //.io_gpio_sws ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561597.4]
  .mem_axi_0_aw_ready ('d1), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_aw_valid (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_aw_bits_id (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_aw_bits_addr (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_aw_bits_len (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_aw_bits_size (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_aw_bits_burst (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_aw_bits_lock (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_aw_bits_cache (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_aw_bits_prot (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_aw_bits_qos (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_w_ready ('d1), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_w_valid (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_w_bits_data (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_w_bits_strb (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_w_bits_last (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_b_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_b_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_b_bits_id ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_b_bits_resp ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_ar_ready ('d1), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_ar_valid (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_ar_bits_id (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_ar_bits_addr (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_ar_bits_len (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_ar_bits_size (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_ar_bits_burst (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_ar_bits_lock (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_ar_bits_cache (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_ar_bits_prot (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_ar_bits_qos (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_r_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_r_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_r_bits_id ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_r_bits_data ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_r_bits_resp ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_0_r_bits_last ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561598.4]
  .mem_axi_1_aw_ready (mem_axi_1_aw_ready), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_aw_valid (mem_axi_1_aw_valid), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_aw_bits_id (mem_axi_1_aw_bits_id), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_aw_bits_addr (mem_axi_1_aw_bits_addr), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_aw_bits_len (mem_axi_1_aw_bits_len), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_aw_bits_size (mem_axi_1_aw_bits_size), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_aw_bits_burst (mem_axi_1_aw_bits_burst), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_aw_bits_lock (mem_axi_1_aw_bits_lock), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_aw_bits_cache (mem_axi_1_aw_bits_cache), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_aw_bits_prot (mem_axi_1_aw_bits_prot), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_aw_bits_qos (mem_axi_1_aw_bits_qos), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_w_ready (mem_axi_1_w_ready), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_w_valid (mem_axi_1_w_valid), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_w_bits_data (mem_axi_1_w_bits_data), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_w_bits_strb (mem_axi_1_w_bits_strb), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_w_bits_last (mem_axi_1_w_bits_last), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_b_ready (mem_axi_1_b_ready), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_b_valid (mem_axi_1_b_valid), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_b_bits_id (mem_axi_1_b_bits_id), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_b_bits_resp (mem_axi_1_b_bits_resp), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_ar_ready (mem_axi_1_ar_ready), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_ar_valid (mem_axi_1_ar_valid), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_ar_bits_id (mem_axi_1_ar_bits_id), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_ar_bits_addr (mem_axi_1_ar_bits_addr), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_ar_bits_len (mem_axi_1_ar_bits_len), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_ar_bits_size (mem_axi_1_ar_bits_size), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_ar_bits_burst (mem_axi_1_ar_bits_burst), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_ar_bits_lock (mem_axi_1_ar_bits_lock), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_ar_bits_cache (mem_axi_1_ar_bits_cache), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_ar_bits_prot (mem_axi_1_ar_bits_prot), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_ar_bits_qos (mem_axi_1_ar_bits_qos), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_r_ready (mem_axi_1_r_ready), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_r_valid (mem_axi_1_r_valid), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_r_bits_id (mem_axi_1_r_bits_id), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_r_bits_data (mem_axi_1_r_bits_data), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_r_bits_resp (mem_axi_1_r_bits_resp), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .mem_axi_1_r_bits_last (mem_axi_1_r_bits_last), // @[:freedom.serve.SERVEiFPGAConfig.fir@561599.4]
  .  mem_axi_2_aw_ready ('d1), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_aw_valid (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_aw_bits_id (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_aw_bits_addr (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_aw_bits_len (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_aw_bits_size (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_aw_bits_burst (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_aw_bits_lock (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_aw_bits_cache (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_aw_bits_prot (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_aw_bits_qos (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_w_ready ('d1), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_w_valid (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_w_bits_data (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_w_bits_strb (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_w_bits_last (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_b_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_b_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_b_bits_id ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_b_bits_resp ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_ar_ready ('d1), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_ar_valid (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_ar_bits_id (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_ar_bits_addr (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_ar_bits_len (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_ar_bits_size (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_ar_bits_burst (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_ar_bits_lock (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_ar_bits_cache (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_ar_bits_prot (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_ar_bits_qos (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_r_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_r_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_r_bits_id ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_r_bits_data ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_r_bits_resp ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mem_axi_2_r_bits_last ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561600.4]
  .mmio_axi_0_aw_ready (mmio_axi_0_aw_ready), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_aw_valid (mmio_axi_0_aw_valid), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_aw_bits_id (mmio_axi_0_aw_bits_id), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_aw_bits_addr (mmio_axi_0_aw_bits_addr), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_aw_bits_len (mmio_axi_0_aw_bits_len), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_aw_bits_size (mmio_axi_0_aw_bits_size), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_aw_bits_burst (mmio_axi_0_aw_bits_burst), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_aw_bits_lock (mmio_axi_0_aw_bits_lock), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_aw_bits_cache (mmio_axi_0_aw_bits_cache), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_aw_bits_prot (mmio_axi_0_aw_bits_prot), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_aw_bits_qos (mmio_axi_0_aw_bits_qos), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_w_ready (mmio_axi_0_w_ready), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_w_valid (mmio_axi_0_w_valid), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_w_bits_data (mmio_axi_0_w_bits_data), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_w_bits_strb (mmio_axi_0_w_bits_strb), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_w_bits_last (mmio_axi_0_w_bits_last), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_b_ready (mmio_axi_0_b_ready), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_b_valid (mmio_axi_0_b_valid), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_b_bits_id (mmio_axi_0_b_bits_id), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_b_bits_resp (mmio_axi_0_b_bits_resp), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_ar_ready (mmio_axi_0_ar_ready), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_ar_valid (mmio_axi_0_ar_valid), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_ar_bits_id (mmio_axi_0_ar_bits_id), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_ar_bits_addr (mmio_axi_0_ar_bits_addr), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_ar_bits_len (mmio_axi_0_ar_bits_len), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_ar_bits_size (mmio_axi_0_ar_bits_size), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_ar_bits_burst (mmio_axi_0_ar_bits_burst), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_ar_bits_lock (mmio_axi_0_ar_bits_lock), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_ar_bits_cache (mmio_axi_0_ar_bits_cache), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_ar_bits_prot (mmio_axi_0_ar_bits_prot), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_ar_bits_qos (mmio_axi_0_ar_bits_qos), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_r_ready (mmio_axi_0_r_ready), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_r_valid (mmio_axi_0_r_valid), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_r_bits_id (mmio_axi_0_r_bits_id), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_r_bits_data (mmio_axi_0_r_bits_data), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_r_bits_resp (mmio_axi_0_r_bits_resp), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  .mmio_axi_0_r_bits_last (mmio_axi_0_r_bits_last), // @[:freedom.serve.SERVEiFPGAConfig.fir@561601.4]
  . front_axi_0_aw_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_aw_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_aw_bits_id ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_aw_bits_addr ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_aw_bits_len ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_aw_bits_size ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_aw_bits_burst ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_aw_bits_lock ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_aw_bits_cache ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_aw_bits_prot ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_aw_bits_qos ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_w_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_w_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_w_bits_data ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_w_bits_strb ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_w_bits_last ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_b_ready ('d1), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_b_valid (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_b_bits_id (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_b_bits_resp (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_ar_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_ar_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_ar_bits_id ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_ar_bits_addr ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_ar_bits_len ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_ar_bits_size ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_ar_bits_burst ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_ar_bits_lock ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_ar_bits_cache ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_ar_bits_prot ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_ar_bits_qos ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_r_ready ('d1), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_r_valid (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_r_bits_id (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_r_bits_data (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_r_bits_resp (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_0_r_bits_last (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561602.4]
  .front_axi_1_aw_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_aw_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_aw_bits_id ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_aw_bits_addr ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_aw_bits_len ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_aw_bits_size ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_aw_bits_burst ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_aw_bits_lock ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_aw_bits_cache ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_aw_bits_prot ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_aw_bits_qos ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_w_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_w_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_w_bits_data ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_w_bits_strb ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_w_bits_last ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_b_ready ('d1), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_b_valid (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_b_bits_id (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_b_bits_resp (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_ar_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_ar_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_ar_bits_id ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_ar_bits_addr ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_ar_bits_len ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_ar_bits_size ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_ar_bits_burst ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_ar_bits_lock ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_ar_bits_cache ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_ar_bits_prot ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_ar_bits_qos ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_r_ready ('d1), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_r_valid (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_r_bits_id (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_r_bits_data (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_r_bits_resp (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_1_r_bits_last (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561603.4]
  .front_axi_2_aw_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_aw_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_aw_bits_id ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_aw_bits_addr ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_aw_bits_len ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_aw_bits_size ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_aw_bits_burst ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_aw_bits_lock ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_aw_bits_cache ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_aw_bits_prot ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_aw_bits_qos ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_w_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_w_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_w_bits_data ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_w_bits_strb ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_w_bits_last ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_b_ready ('d1), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_b_valid (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_b_bits_id (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_b_bits_resp (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_ar_ready (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_ar_valid ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_ar_bits_id ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_ar_bits_addr ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_ar_bits_len ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_ar_bits_size ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_ar_bits_burst ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_ar_bits_lock ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_ar_bits_cache ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_ar_bits_prot ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_ar_bits_qos ('d0), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_r_ready ('d1), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_r_valid (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_r_bits_id (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_r_bits_data (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_r_bits_resp (), // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
  .front_axi_2_r_bits_last () // @[:freedom.serve.SERVEiFPGAConfig.fir@561604.4]
);
endmodule